module mux31x64 (dataout, a, b, c, s);

   input [63:0]  a, b, c;
   input [1:0] 	 s;

   output [63:0] dataout;

   mux31 m1 (dataout[0], a[0], b[0], c[0], s);
   mux31 m2 (dataout[1], a[1], b[1], c[1], s);
   mux31 m3 (dataout[2], a[2], b[2], c[2], s);
   mux31 m4 (dataout[3], a[3], b[3], c[3], s);
   mux31 m5 (dataout[4], a[4], b[4], c[4], s);
   mux31 m6 (dataout[5], a[5], b[5], c[5], s);
   mux31 m7 (dataout[6], a[6], b[6], c[6], s);
   mux31 m8 (dataout[7], a[7], b[7], c[7], s);
   mux31 m9 (dataout[8], a[8], b[8], c[8], s);
   mux31 m10 (dataout[9], a[9], b[9], c[9], s);
   mux31 m11 (dataout[10], a[10], b[10], c[10], s);
   mux31 m12 (dataout[11], a[11], b[11], c[11], s);
   mux31 m13 (dataout[12], a[12], b[12], c[12], s);
   mux31 m14 (dataout[13], a[13], b[13], c[13], s);
   mux31 m15 (dataout[14], a[14], b[14], c[14], s);
   mux31 m16 (dataout[15], a[15], b[15], c[15], s);
   mux31 m17 (dataout[16], a[16], b[16], c[16], s);
   mux31 m18 (dataout[17], a[17], b[17], c[17], s);
   mux31 m19 (dataout[18], a[18], b[18], c[18], s);
   mux31 m20 (dataout[19], a[19], b[19], c[19], s);
   mux31 m21 (dataout[20], a[20], b[20], c[20], s);
   mux31 m22 (dataout[21], a[21], b[21], c[21], s);
   mux31 m23 (dataout[22], a[22], b[22], c[22], s);
   mux31 m24 (dataout[23], a[23], b[23], c[23], s);
   mux31 m25 (dataout[24], a[24], b[24], c[24], s);
   mux31 m26 (dataout[25], a[25], b[25], c[25], s);
   mux31 m27 (dataout[26], a[26], b[26], c[26], s);
   mux31 m28 (dataout[27], a[27], b[27], c[27], s);
   mux31 m29 (dataout[28], a[28], b[28], c[28], s);
   mux31 m30 (dataout[29], a[29], b[29], c[29], s);
   mux31 m31 (dataout[30], a[30], b[30], c[30], s);
   mux31 m32 (dataout[31], a[31], b[31], c[31], s);
   mux31 m33 (dataout[32], a[32], b[32], c[32], s);
   mux31 m34 (dataout[33], a[33], b[33], c[33], s);
   mux31 m35 (dataout[34], a[34], b[34], c[34], s);
   mux31 m36 (dataout[35], a[35], b[35], c[35], s);
   mux31 m37 (dataout[36], a[36], b[36], c[36], s);
   mux31 m38 (dataout[37], a[37], b[37], c[37], s);
   mux31 m39 (dataout[38], a[38], b[38], c[38], s);
   mux31 m40 (dataout[39], a[39], b[39], c[39], s);
   mux31 m41 (dataout[40], a[40], b[40], c[40], s);
   mux31 m42 (dataout[41], a[41], b[41], c[41], s);
   mux31 m43 (dataout[42], a[42], b[42], c[42], s);
   mux31 m44 (dataout[43], a[43], b[43], c[43], s);
   mux31 m45 (dataout[44], a[44], b[44], c[44], s);
   mux31 m46 (dataout[45], a[45], b[45], c[45], s);
   mux31 m47 (dataout[46], a[46], b[46], c[46], s);
   mux31 m48 (dataout[47], a[47], b[47], c[47], s);
   mux31 m49 (dataout[48], a[48], b[48], c[48], s);
   mux31 m50 (dataout[49], a[49], b[49], c[49], s);
   mux31 m51 (dataout[50], a[50], b[50], c[50], s);
   mux31 m52 (dataout[51], a[51], b[51], c[51], s);
   mux31 m53 (dataout[52], a[52], b[52], c[52], s);
   mux31 m54 (dataout[53], a[53], b[53], c[53], s);
   mux31 m55 (dataout[54], a[54], b[54], c[54], s);
   mux31 m56 (dataout[55], a[55], b[55], c[55], s);
   mux31 m57 (dataout[56], a[56], b[56], c[56], s);
   mux31 m58 (dataout[57], a[57], b[57], c[57], s);
   mux31 m59 (dataout[58], a[58], b[58], c[58], s);
   mux31 m60 (dataout[59], a[59], b[59], c[59], s);
   mux31 m61 (dataout[60], a[60], b[60], c[60], s);
   mux31 m62 (dataout[61], a[61], b[61], c[61], s);
   mux31 m63 (dataout[62], a[62], b[62], c[62], s);
   mux31 m64 (dataout[63], a[63], b[63], c[63], s);

endmodule // mux31x64
